
module unsaved (
	clk_clk,
	reset_reset_n,
	leds_out_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[9:0]	leds_out_export;
endmodule
